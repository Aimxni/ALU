module shifter(in,shift,sout);
input [15:0] in;
input [1:0] shift;
output [15:0] sout;
reg [15:0] sout;



// fill outhe rest
always_comb 
begin 
    
    if (shift == 2'b00)
        sout = in;
    else if (shift == 2'b01)
        sout = in << 1;
    else if (shift == 2'b10)
        sout = in >> 1;
    else if (shift == 2'b11)
    begin
      sout = in >> 1;
      sout[15] = in[15];
    end 
    else 
    sout = 16'bxxxxxxxxxxxxxxxx;




end 
endmodule